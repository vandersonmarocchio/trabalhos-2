CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
55
13 Logic Switch~
5 693 127 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8152 0 0
2
5.89895e-315 0
0
13 Logic Switch~
5 663 127 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 Cin
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6223 0 0
2
5.89895e-315 0
0
13 Logic Switch~
5 724 126 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5441 0 0
2
5.89895e-315 0
0
13 Logic Switch~
5 235 130 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3189 0 0
2
5.89895e-315 5.30499e-315
0
13 Logic Switch~
5 299 129 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8460 0 0
2
5.89895e-315 5.26354e-315
0
13 Logic Switch~
5 361 130 0 10 11
0 52 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5179 0 0
2
5.89895e-315 0
0
9 Inverter~
13 690 751 0 2 22
0 7 6
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3593 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 975 786 0 3 22
0 12 2 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SUB
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
3928 0 0
2
5.89895e-315 5.37752e-315
0
9 2-In AND~
219 973 865 0 3 22
0 2 13 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SUB
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
363 0 0
2
5.89895e-315 5.36716e-315
0
8 3-In OR~
219 868 874 0 4 22
0 10 11 9 13
0
0 0 624 0
4 4075
-14 -24 14 -16
3 SUB
-1 -4 20 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 13 0
1 U
8132 0 0
2
5.89895e-315 5.3568e-315
0
9 2-In AND~
219 765 914 0 3 22
0 8 6 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SUB
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
65 0 0
2
5.89895e-315 5.34643e-315
0
9 2-In AND~
219 765 875 0 3 22
0 6 5 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SUB
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
6609 0 0
2
5.89895e-315 5.32571e-315
0
9 2-In AND~
219 765 833 0 3 22
0 8 5 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SUB
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
8995 0 0
2
5.89895e-315 5.30499e-315
0
6 74136~
219 869 777 0 3 22
0 7 14 12
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUB
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
3918 0 0
2
5.89895e-315 5.26354e-315
0
6 74136~
219 758 787 0 3 22
0 8 5 14
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SUB
-2 -5 19 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
7519 0 0
2
5.89895e-315 0
0
14 Logic Display~
6 1121 707 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
4 Cout
-13 -26 15 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
377 0 0
2
5.89895e-315 0
0
14 Logic Display~
6 1122 637 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 S
-3 -26 4 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8816 0 0
2
5.89895e-315 0
0
8 2-In OR~
219 1063 732 0 3 22
0 17 3 16
0
0 0 112 0
6 74LS32
-21 -24 21 -16
2 A1
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
3877 0 0
2
5.89895e-315 0
0
8 2-In OR~
219 1063 655 0 3 22
0 18 4 15
0
0 0 112 0
6 74LS32
-21 -24 21 -16
2 A2
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
926 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 975 522 0 3 22
0 23 19 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SOM
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
7262 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 973 601 0 3 22
0 19 24 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SOM
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
5267 0 0
2
5.89895e-315 0
0
8 3-In OR~
219 868 610 0 4 22
0 21 22 20 24
0
0 0 624 0
4 4075
-14 -24 14 -16
3 SOM
-1 -4 20 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 13 0
1 U
8838 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 765 650 0 3 22
0 8 7 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SOM
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
7159 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 765 611 0 3 22
0 7 5 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SOM
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
5812 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 765 569 0 3 22
0 8 5 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 SOM
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
331 0 0
2
5.89895e-315 0
0
6 74136~
219 869 513 0 3 22
0 7 25 23
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SOM
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
9604 0 0
2
5.89895e-315 0
0
6 74136~
219 758 523 0 3 22
0 8 5 25
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 SOM
-2 -5 19 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
7518 0 0
2
5.89895e-315 0
0
14 Logic Display~
6 1112 303 0 1 2
10 34
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 R3
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4832 0 0
2
5.89895e-315 0
0
8 3-In OR~
219 1043 326 0 4 22
0 27 35 26 34
0
0 0 112 0
4 4075
-14 -24 14 -16
2 A4
-7 -34 7 -26
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 13 0
1 U
6798 0 0
2
5.89895e-315 0
0
8 2-In OR~
219 916 415 0 3 22
0 29 28 26
0
0 0 112 0
6 74LS32
-21 -24 21 -16
2 A5
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3336 0 0
2
5.89895e-315 0
0
8 2-In OR~
219 919 325 0 3 22
0 31 30 35
0
0 0 112 0
6 74LS32
-21 -24 21 -16
2 A6
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
8370 0 0
2
5.89895e-315 0
0
8 2-In OR~
219 918 245 0 3 22
0 33 32 27
0
0 0 112 0
6 74LS32
-21 -24 21 -16
2 A7
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3910 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 759 216 0 3 22
0 7 5 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
316 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 828 395 0 3 22
0 42 37 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 XOR
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
536 0 0
2
5.89895e-315 5.36716e-315
0
9 2-In AND~
219 830 440 0 3 22
0 41 36 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 XNOR
-17 -2 11 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
4460 0 0
2
5.89895e-315 5.3568e-315
0
9 2-In AND~
219 828 304 0 3 22
0 44 39 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 OR
-10 -4 4 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3260 0 0
2
5.89895e-315 5.30499e-315
0
9 2-In AND~
219 828 347 0 3 22
0 43 38 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 NOR
-14 -3 7 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5156 0 0
2
5.89895e-315 5.26354e-315
0
9 2-In AND~
219 829 263 0 3 22
0 45 40 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 NAND
-17 -3 11 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3133 0 0
2
5.89895e-315 0
0
9 2-In AND~
219 828 225 0 3 22
0 46 47 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
5523 0 0
2
5.89895e-315 5.37752e-315
0
6 74266~
219 752 431 0 3 22
0 7 5 41
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 XNOR
-3 -4 25 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3746 0 0
2
5.89895e-315 5.34643e-315
0
6 74136~
219 751 386 0 3 22
0 7 5 42
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 XOR
-1 -5 20 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
5668 0 0
2
5.89895e-315 5.32571e-315
0
9 2-In NOR~
219 748 338 0 3 22
0 7 5 43
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 NOR
-2 -4 19 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
5368 0 0
2
5.89895e-315 5.30499e-315
0
8 2-In OR~
219 749 295 0 3 22
0 7 5 44
0
0 0 624 0
6 74LS32
-21 -24 21 -16
2 OR
1 -4 15 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8293 0 0
2
5.89895e-315 5.26354e-315
0
10 2-In NAND~
219 758 254 0 3 22
0 7 5 45
0
0 0 624 0
4 7400
-7 -24 21 -16
4 NAND
-16 -4 12 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3232 0 0
2
5.89895e-315 0
0
9 Inverter~
13 257 181 0 2 22
0 48 49
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6644 0 0
2
5.89895e-315 5.41378e-315
0
9 Inverter~
13 321 180 0 2 22
0 50 51
0
0 0 112 270
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4978 0 0
2
5.89895e-315 5.4086e-315
0
9 Inverter~
13 383 181 0 2 22
0 52 53
0
0 0 112 270
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9207 0 0
2
5.89895e-315 5.40342e-315
0
5 7415~
219 434 216 0 4 22
0 49 51 53 47
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 AND
-13 -4 8 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
6998 0 0
2
5.89895e-315 5.39824e-315
0
5 7415~
219 435 257 0 4 22
0 49 51 52 40
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 NAND
-16 -2 12 6
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
3175 0 0
2
5.89895e-315 5.39306e-315
0
5 7415~
219 435 298 0 4 22
0 49 50 53 39
0
0 0 624 0
6 74LS15
-21 -28 21 -20
2 OR
-10 -3 4 5
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
3378 0 0
2
5.89895e-315 5.38788e-315
0
5 7415~
219 435 341 0 4 22
0 49 50 52 38
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 NOR
-13 -3 8 5
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
922 0 0
2
5.89895e-315 5.37752e-315
0
5 7415~
219 432 527 0 4 22
0 48 50 52 2
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 SUB
-13 -3 8 5
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
6891 0 0
2
5.89895e-315 5.36716e-315
0
5 7415~
219 433 481 0 4 22
0 48 50 53 19
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 SOM
-13 -4 8 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 3 0
1 U
5407 0 0
2
5.89895e-315 5.3568e-315
0
5 7415~
219 434 434 0 4 22
0 48 51 52 36
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 XNOR
-15 -5 13 3
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
7349 0 0
2
5.89895e-315 5.34643e-315
0
5 7415~
219 435 389 0 4 22
0 48 51 53 37
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 XOR
-12 -4 9 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 4 0
1 U
3919 0 0
2
5.89895e-315 5.32571e-315
0
111
1 0 2 0 0 8192 0 9 0 0 4 3
949 856
900 856
900 795
3 2 3 0 0 8320 0 9 18 0 0 4
994 865
1027 865
1027 741
1050 741
3 2 4 0 0 8320 0 8 19 0 0 4
996 786
1013 786
1013 664
1050 664
2 4 2 0 0 12416 0 8 52 0 0 6
951 795
791 795
791 811
481 811
481 527
453 527
2 0 5 0 0 4096 0 12 0 0 17 2
741 884
724 884
2 0 5 0 0 0 0 13 0 0 17 2
741 842
724 842
2 0 5 0 0 4096 0 15 0 0 17 2
742 796
724 796
2 0 5 0 0 0 0 24 0 0 17 2
741 620
724 620
2 0 5 0 0 0 0 25 0 0 17 2
741 578
724 578
2 0 5 0 0 0 0 27 0 0 17 2
742 532
724 532
2 0 5 0 0 0 0 40 0 0 17 2
736 440
724 440
2 0 5 0 0 0 0 41 0 0 17 2
735 395
724 395
2 0 5 0 0 0 0 42 0 0 17 2
735 347
724 347
2 0 5 0 0 0 0 43 0 0 17 2
736 304
724 304
2 0 5 0 0 0 0 44 0 0 17 2
734 263
724 263
2 0 5 0 0 0 0 33 0 0 17 2
735 225
724 225
1 0 5 0 0 4224 0 3 0 0 0 2
724 138
724 952
2 0 6 0 0 4096 0 11 0 0 30 2
741 923
693 923
1 0 6 0 0 0 0 12 0 0 30 2
741 866
693 866
1 0 7 0 0 12288 0 14 0 0 31 4
853 768
806 768
806 717
693 717
2 0 7 0 0 0 0 23 0 0 31 2
741 659
693 659
1 0 7 0 0 0 0 24 0 0 31 2
741 602
693 602
1 0 7 0 0 0 0 26 0 0 31 4
853 504
805 504
805 475
693 475
1 0 7 0 0 0 0 40 0 0 31 2
736 422
693 422
1 0 7 0 0 0 0 41 0 0 31 2
735 377
693 377
1 0 7 0 0 0 0 42 0 0 31 2
735 329
693 329
1 0 7 0 0 0 0 43 0 0 31 2
736 286
693 286
1 0 7 0 0 0 0 44 0 0 31 2
734 245
693 245
1 0 7 0 0 0 0 33 0 0 31 2
735 207
693 207
2 0 6 0 0 4224 0 7 0 0 0 2
693 769
693 951
1 1 7 0 0 4224 0 1 7 0 0 2
693 139
693 733
1 0 8 0 0 4096 0 11 0 0 38 2
741 905
663 905
1 0 8 0 0 0 0 13 0 0 38 2
741 824
663 824
1 0 8 0 0 4096 0 15 0 0 38 2
742 778
663 778
1 0 8 0 0 0 0 23 0 0 38 2
741 641
663 641
1 0 8 0 0 0 0 25 0 0 38 2
741 560
663 560
1 0 8 0 0 0 0 27 0 0 38 2
742 514
663 514
1 0 8 0 0 4224 0 2 0 0 0 2
663 139
663 953
3 3 9 0 0 4224 0 10 11 0 0 4
855 883
806 883
806 914
786 914
3 1 10 0 0 12416 0 13 10 0 0 4
786 833
806 833
806 865
855 865
2 3 11 0 0 4224 0 10 12 0 0 3
856 874
786 874
786 875
1 3 12 0 0 4224 0 8 14 0 0 2
951 777
902 777
2 4 13 0 0 4224 0 9 10 0 0 2
949 874
901 874
2 3 14 0 0 4224 0 14 15 0 0 3
853 786
791 786
791 787
1 3 15 0 0 4224 0 17 19 0 0 2
1122 655
1096 655
1 3 16 0 0 8320 0 16 18 0 0 3
1121 725
1121 732
1096 732
3 1 17 0 0 8320 0 21 18 0 0 4
994 601
1001 601
1001 723
1050 723
3 1 18 0 0 8320 0 20 19 0 0 4
996 522
1028 522
1028 646
1050 646
1 0 19 0 0 8192 0 21 0 0 53 3
949 592
900 592
900 531
3 3 20 0 0 4224 0 22 23 0 0 4
855 619
806 619
806 650
786 650
3 1 21 0 0 12416 0 25 22 0 0 4
786 569
806 569
806 601
855 601
2 3 22 0 0 4224 0 22 24 0 0 3
856 610
786 610
786 611
2 4 19 0 0 12416 0 20 53 0 0 6
951 531
791 531
791 546
512 546
512 481
454 481
1 3 23 0 0 4224 0 20 26 0 0 2
951 513
902 513
2 4 24 0 0 4224 0 21 22 0 0 2
949 610
901 610
2 3 25 0 0 4224 0 26 27 0 0 3
853 522
791 522
791 523
3 3 26 0 0 8320 0 29 30 0 0 4
1030 335
997 335
997 415
949 415
1 3 27 0 0 8320 0 29 32 0 0 4
1030 317
997 317
997 245
951 245
3 2 28 0 0 12416 0 35 30 0 0 4
851 440
875 440
875 424
903 424
1 3 29 0 0 4224 0 30 34 0 0 4
903 406
875 406
875 395
849 395
3 2 30 0 0 12416 0 37 31 0 0 4
849 347
875 347
875 334
906 334
3 1 31 0 0 12416 0 36 31 0 0 4
849 304
875 304
875 316
906 316
2 3 32 0 0 4224 0 32 38 0 0 4
905 254
875 254
875 263
850 263
3 1 33 0 0 12416 0 39 32 0 0 4
849 225
875 225
875 236
905 236
1 4 34 0 0 8320 0 28 29 0 0 3
1112 321
1112 326
1076 326
2 3 35 0 0 4224 0 29 31 0 0 4
1031 326
967 326
967 325
952 325
4 2 36 0 0 12416 0 54 35 0 0 4
455 434
530 434
530 449
806 449
2 4 37 0 0 4224 0 34 55 0 0 4
804 404
554 404
554 389
456 389
2 4 38 0 0 4224 0 37 51 0 0 4
804 356
584 356
584 341
456 341
2 4 39 0 0 4224 0 36 50 0 0 4
804 313
598 313
598 298
456 298
2 4 40 0 0 4224 0 38 49 0 0 4
805 272
618 272
618 257
456 257
3 1 41 0 0 4224 0 40 35 0 0 2
791 431
806 431
3 1 42 0 0 4224 0 41 34 0 0 2
784 386
804 386
3 1 43 0 0 4224 0 42 37 0 0 2
787 338
804 338
3 1 44 0 0 4224 0 43 36 0 0 2
782 295
804 295
3 1 45 0 0 4224 0 44 38 0 0 2
785 254
805 254
3 1 46 0 0 4224 0 33 39 0 0 2
780 216
804 216
4 2 47 0 0 4224 0 48 39 0 0 4
455 216
636 216
636 234
804 234
1 0 48 0 0 4096 0 52 0 0 111 2
408 518
235 518
1 0 48 0 0 4096 0 53 0 0 111 2
409 472
235 472
1 0 48 0 0 4096 0 54 0 0 111 2
410 425
235 425
1 0 48 0 0 4096 0 55 0 0 111 2
411 380
235 380
1 0 49 0 0 4096 0 51 0 0 109 2
411 332
260 332
1 0 49 0 0 0 0 50 0 0 109 2
411 289
260 289
1 0 49 0 0 0 0 49 0 0 109 2
411 248
260 248
2 0 50 0 0 4096 0 52 0 0 108 2
408 527
299 527
2 0 50 0 0 4096 0 53 0 0 108 2
409 481
299 481
2 0 51 0 0 4096 0 54 0 0 106 2
410 434
324 434
2 0 51 0 0 4096 0 55 0 0 106 2
411 389
324 389
2 0 50 0 0 4096 0 51 0 0 108 2
411 341
299 341
2 0 50 0 0 0 0 50 0 0 108 2
411 298
299 298
2 0 51 0 0 0 0 49 0 0 106 2
411 257
324 257
3 0 52 0 0 4096 0 52 0 0 105 2
408 536
361 536
3 0 53 0 0 4096 0 53 0 0 103 2
409 490
386 490
3 0 52 0 0 4096 0 54 0 0 105 2
410 443
361 443
3 0 53 0 0 4096 0 55 0 0 103 2
411 398
386 398
3 0 52 0 0 4096 0 51 0 0 105 2
411 350
361 350
3 0 53 0 0 0 0 50 0 0 103 2
411 307
386 307
3 0 52 0 0 0 0 49 0 0 105 2
411 266
361 266
3 0 53 0 0 0 0 48 0 0 103 2
410 225
386 225
2 0 51 0 0 0 0 48 0 0 106 2
410 216
324 216
1 0 49 0 0 0 0 48 0 0 109 2
410 207
260 207
2 0 53 0 0 4224 0 47 0 0 0 2
386 199
386 556
1 0 52 0 0 0 0 47 0 0 105 2
386 163
361 163
1 0 52 0 0 4224 0 6 0 0 0 2
361 142
361 556
2 0 51 0 0 4224 0 46 0 0 0 2
324 198
324 555
1 0 50 0 0 0 0 46 0 0 108 2
324 162
299 162
1 0 50 0 0 4224 0 5 0 0 0 2
299 141
299 555
2 0 49 0 0 4224 0 45 0 0 0 2
260 199
260 556
1 0 48 0 0 0 0 45 0 0 111 2
260 163
235 163
1 0 48 0 0 4224 0 4 0 0 0 2
235 142
235 556
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 95
108 203 217 387
118 211 206 355
95 000 -> AND
001 -> NAND
010 -> OR
011 -> NOR
100 -> XOR
101 -> XNOR
110 -> SOM
111 -> SUB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1065 260 1182 284
1075 268 1171 284
12 Sa�da L�gica
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
651 59 736 83
661 67 725 83
8 Entradas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
244 62 369 86
254 70 358 86
13 Decocificador
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
731 161 872 185
741 169 861 185
15 Fun��es L�gicas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1058 575 1207 599
1068 583 1196 599
16 Sa�da Aritm�tica
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
