CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
37
13 Logic Switch~
5 311 551 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 CS
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89906e-315 5.3568e-315
0
13 Logic Switch~
5 312 588 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 RD
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89906e-315 5.34643e-315
0
13 Logic Switch~
5 311 628 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 OE
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89906e-315 5.32571e-315
0
13 Logic Switch~
5 310 296 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89906e-315 0
0
13 Logic Switch~
5 625 228 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 E0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89906e-315 5.34643e-315
0
13 Logic Switch~
5 755 234 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 E1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89906e-315 5.32571e-315
0
13 Logic Switch~
5 887 229 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 E2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.89906e-315 5.30499e-315
0
9 Inverter~
13 406 474 0 2 22
0 4 5
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 2 0
1 U
7361 0 0
2
5.89906e-315 0
0
12 D Flip-Flop~
219 941 437 0 4 9
0 33 32 36 6
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.89906e-315 0
0
12 D Flip-Flop~
219 798 435 0 4 9
0 34 32 37 8
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U5
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
972 0 0
2
5.89906e-315 0
0
12 D Flip-Flop~
219 673 432 0 4 9
0 35 32 38 10
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U4
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89906e-315 0
0
12 D Flip-Flop~
219 935 355 0 4 9
0 33 31 39 7
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
5.89906e-315 0
0
12 D Flip-Flop~
219 803 356 0 4 9
0 34 31 40 9
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.89906e-315 0
0
12 D Flip-Flop~
219 675 355 0 4 9
0 35 31 41 11
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4597 0 0
2
5.89906e-315 0
0
9 Inverter~
13 390 242 0 2 22
0 13 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 2 0
1 U
3835 0 0
2
5.89906e-315 0
0
14 Logic Display~
6 1396 246 0 1 2
31 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 D0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.89906e-315 5.41896e-315
0
9 2-In AND~
219 1182 260 0 3 22
0 11 12 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 CC
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
5616 0 0
2
5.89906e-315 5.41378e-315
0
9 2-In AND~
219 1183 308 0 3 22
0 10 13 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 CD
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9323 0 0
2
5.89906e-315 5.4086e-315
0
9 2-In AND~
219 1185 432 0 3 22
0 8 13 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 C1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
317 0 0
2
5.89906e-315 5.40342e-315
0
9 2-In AND~
219 1184 384 0 3 22
0 9 12 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 C1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3108 0 0
2
5.89906e-315 5.39824e-315
0
9 2-In AND~
219 1186 563 0 3 22
0 6 13 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 C1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
4299 0 0
2
5.89906e-315 5.39306e-315
0
9 2-In AND~
219 1185 515 0 3 22
0 7 12 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 C1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9672 0 0
2
5.89906e-315 5.38788e-315
0
8 2-In OR~
219 1258 269 0 3 22
0 27 26 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7876 0 0
2
5.89906e-315 5.37752e-315
0
8 2-In OR~
219 1264 393 0 3 22
0 25 23 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
6369 0 0
2
5.89906e-315 5.36716e-315
0
8 2-In OR~
219 1266 524 0 3 22
0 24 22 19
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9172 0 0
2
5.89906e-315 5.3568e-315
0
10 Buffer 3S~
219 1326 269 0 3 22
0 21 15 18
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
6 BuffeB
-21 -20 21 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7100 0 0
2
5.89906e-315 5.34643e-315
0
10 Buffer 3S~
219 1333 393 0 3 22
0 20 15 17
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
6 BuffeC
-21 -20 21 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3820 0 0
2
5.89906e-315 5.32571e-315
0
10 Buffer 3S~
219 1338 524 0 3 22
0 19 15 16
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
6 BuffeD
-21 -20 21 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
7678 0 0
2
5.89906e-315 5.30499e-315
0
14 Logic Display~
6 1402 370 0 1 2
31 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 D1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89906e-315 5.26354e-315
0
14 Logic Display~
6 1408 501 0 1 2
31 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 D2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.89906e-315 0
0
9 Inverter~
13 356 551 0 2 22
0 30 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3409 0 0
2
5.89906e-315 5.30499e-315
0
9 Inverter~
13 381 627 0 2 22
0 29 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 2 0
1 U
3951 0 0
2
5.89906e-315 5.26354e-315
0
5 7415~
219 497 560 0 4 22
0 14 4 28 15
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
8885 0 0
2
5.89906e-315 0
0
9 2-In AND~
219 533 250 0 3 22
0 12 2 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 CC
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3780 0 0
2
5.89906e-315 5.26354e-315
0
9 2-In AND~
219 534 304 0 3 22
0 13 2 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 CB
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9265 0 0
2
5.89906e-315 0
0
7 Pulser~
4 330 349 0 10 12
0 42 43 44 3 0 0 10 10 10
7
0
0 0 4656 0
0
6 Pulser
-21 -28 21 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9442 0 0
2
5.89906e-315 5.40342e-315
0
5 7415~
219 463 396 0 4 22
0 3 14 5 2
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
9424 0 0
2
5.89906e-315 5.34643e-315
0
53
2 0 2 0 0 4096 0 35 0 0 2 2
510 313
498 313
4 2 2 0 0 8320 0 37 34 0 0 4
484 396
498 396
498 259
509 259
4 1 3 0 0 4224 0 36 37 0 0 4
360 349
420 349
420 387
439 387
1 0 4 0 0 4096 0 8 0 0 37 3
409 492
409 560
408 560
2 3 5 0 0 4224 0 8 37 0 0 3
409 456
409 405
439 405
4 1 6 0 0 8320 0 9 21 0 0 6
965 401
992 401
992 626
1078 626
1078 554
1162 554
4 1 7 0 0 8320 0 12 22 0 0 6
959 319
982 319
982 636
1087 636
1087 506
1161 506
4 1 8 0 0 20608 0 10 19 0 0 6
822 399
860 399
860 517
1009 517
1009 423
1161 423
4 1 9 0 0 8320 0 13 20 0 0 6
827 320
844 320
844 528
1019 528
1019 375
1160 375
4 1 10 0 0 12416 0 11 18 0 0 6
697 396
729 396
729 551
1048 551
1048 299
1159 299
4 1 11 0 0 12416 0 14 17 0 0 6
699 319
716 319
716 562
1061 562
1061 251
1158 251
2 0 12 0 0 4096 0 20 0 0 17 2
1160 393
1107 393
2 0 12 0 0 0 0 17 0 0 17 2
1158 269
1107 269
2 0 13 0 0 4096 0 18 0 0 16 2
1159 317
1143 317
2 0 13 0 0 4096 0 19 0 0 16 2
1161 441
1143 441
0 2 13 0 0 8320 0 0 21 41 0 5
332 296
332 155
1143 155
1143 572
1162 572
0 2 12 0 0 8320 0 0 22 19 0 5
417 242
417 165
1107 165
1107 524
1161 524
1 0 13 0 0 0 0 15 0 0 41 3
375 242
347 242
347 296
2 1 12 0 0 0 0 15 34 0 0 4
411 242
417 242
417 241
509 241
2 0 14 0 0 8320 0 37 0 0 38 3
439 396
390 396
390 551
2 0 15 0 0 8192 0 28 0 0 23 3
1338 535
1338 579
1440 579
2 0 15 0 0 8192 0 27 0 0 23 3
1333 404
1333 446
1440 446
4 2 15 0 0 12416 0 33 26 0 0 7
518 560
705 560
705 648
1440 648
1440 293
1326 293
1326 280
1 3 16 0 0 8320 0 30 28 0 0 3
1408 519
1408 524
1353 524
1 3 17 0 0 8320 0 29 27 0 0 3
1402 388
1402 393
1348 393
1 3 18 0 0 8320 0 16 26 0 0 3
1396 264
1396 269
1341 269
1 3 19 0 0 4224 0 28 25 0 0 2
1323 524
1299 524
3 1 20 0 0 4224 0 24 27 0 0 2
1297 393
1318 393
1 3 21 0 0 4224 0 26 23 0 0 2
1311 269
1291 269
3 2 22 0 0 8320 0 21 25 0 0 4
1207 563
1233 563
1233 533
1253 533
3 2 23 0 0 8320 0 19 24 0 0 4
1206 432
1233 432
1233 402
1251 402
1 3 24 0 0 4224 0 25 22 0 0 2
1253 515
1206 515
1 3 25 0 0 4224 0 24 20 0 0 2
1251 384
1205 384
3 2 26 0 0 8320 0 18 23 0 0 4
1204 308
1232 308
1232 278
1245 278
3 1 27 0 0 4224 0 17 23 0 0 2
1203 260
1245 260
2 3 28 0 0 8320 0 32 33 0 0 4
402 627
440 627
440 569
473 569
1 2 4 0 0 4224 0 2 33 0 0 4
324 588
408 588
408 560
473 560
1 2 14 0 0 0 0 33 31 0 0 2
473 551
377 551
1 1 29 0 0 8320 0 3 32 0 0 3
323 628
323 627
366 627
1 1 30 0 0 4224 0 31 1 0 0 4
341 551
322 551
322 551
323 551
1 1 13 0 0 0 0 35 4 0 0 4
510 295
347 295
347 296
322 296
2 0 31 0 0 8192 0 14 0 0 44 3
651 337
607 337
607 251
2 0 31 0 0 8192 0 13 0 0 44 3
779 338
739 338
739 251
3 2 31 0 0 12416 0 34 12 0 0 6
554 250
607 250
607 251
872 251
872 337
911 337
2 0 32 0 0 8192 0 11 0 0 47 3
649 414
602 414
602 491
2 0 32 0 0 0 0 10 0 0 47 3
774 417
740 417
740 491
3 2 32 0 0 12416 0 35 9 0 0 6
555 304
563 304
563 491
887 491
887 419
917 419
1 0 33 0 0 4096 0 12 0 0 49 2
911 319
888 319
1 1 33 0 0 12416 0 7 9 0 0 5
887 241
887 319
888 319
888 401
917 401
1 0 34 0 0 4096 0 13 0 0 51 2
779 320
755 320
1 1 34 0 0 4224 0 6 10 0 0 3
755 246
755 399
774 399
1 0 35 0 0 4096 0 14 0 0 53 2
651 319
626 319
1 1 35 0 0 4224 0 5 11 0 0 5
625 240
625 319
626 319
626 396
649 396
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
228 222 305 246
238 230 294 246
7 ENTRADA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
217 237 326 261
227 245 315 261
11 DE ENDERE�O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
210 491 367 515
220 499 356 515
17 LEITURA E ESCRITA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
232 476 341 500
242 484 330 500
11 CONTROLE DE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
688 168 837 192
698 176 826 192
16 LEITURA DE DADOS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1229 194 1306 218
1239 202 1295 218
7 ESCRITA
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
